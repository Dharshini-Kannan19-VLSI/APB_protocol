 package APB_Pkg;
    import uvm_pkg::*;
   `include "uvm_macros.svh"

 //Include all files
   `include "APB_Transaction.sv"
   `include "APB_Sequence.sv"
   `include "APB_Sequencer.sv"
   `include "APB_Driver.sv"
   `include "APB_Monitor.sv"
   `include "APB_Agent.sv"
   `include "APB_Scoreboard.sv"
   `include "APB_Env.sv"
   `include "APB_Test.sv"
endpackage